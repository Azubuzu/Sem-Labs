--
-- VHDL Architecture Morse.charToMorseController.studentVersion
--
-- Created:
--          by - leo.dosreis.UNKNOWN (WE5400)
--          at - 11:19:15 25.04.2018
--
-- using Mentor Graphics HDL Designer(TM) 2015.2 (Build 5)
--
ARCHITECTURE studentVersion OF charToMorseController IS
BEGIN
END ARCHITECTURE studentVersion;

